module top;
	/**************************** TIMING DECLARATION ******************************/
    timeunit 1ns;
    timeprecision 1ns;
    int timeout = 1000000;

    /***************************** CLOCK GENERATION *******************************/
    bit clk;
    always #5 clk = clk === 1'b0;

    /*************************** TESTBENCH DECLARATION ****************************/
    two_bit_multiplier_tb tb_i(.*);

	/******************************* TIME OUT TRAP ********************************/
    always @(posedge clk) begin
		if (timeout == 0) begin
			// $display("		Timed out ⏳⏳⏳ ❌ ❌ ❌");
			// $finish;
		end
		timeout <= timeout - 1;
	end

	/**************************** INITIAL DECLARATION ******************************/
    initial begin
		$dumpfile("waveform.vcd");
		$dumpvars();

		tb_i.main();

		$display("		SUCCESS!!! 💯 💯 💯 ✅ ✅ ✅");
		$finish;
	end

endmodule